`ifndef __INCLUDE_VH__
`define __INCLUDE_VH__

`include "./headers/ISA.svh"
`include "./headers/sys_defs.svh"
`include "./headers/fetch_defs.svh"
`include "./headers/execute.svh"
`include "./headers/dispatch_defs.svh"
`include "./headers/issue_defs.svh"
`include "./headers/pipeline_defs.svh"

`endif
